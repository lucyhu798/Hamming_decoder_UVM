// Code your testbench here
// or browse Examples
`define QUESTA
`include "hamming_pkg.sv"
`include "hamming_bfm.sv"
`include "top.sv"
