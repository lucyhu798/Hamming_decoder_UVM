/*
   Copyright 2013 Ray Salemi
*/
package hamming_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
`include "transaction.sv"
`include "coverage.sv"
`include "scoreboard.sv"
`include "result_monitor.sv"
`include "h_sequencer.sv"
`include "driver.sv"
`include "hamming_agent.sv"
`include "env.sv"
`include "no_error_sequence.sv"
`include "one_error_sequence.sv"
`include "two_error_sequence.sv"
`include "no_error_test.sv"
`include "one_error_test.sv"
`include "two_error_test.sv"
   
endpackage : hamming_pkg

   